// testbench for gpsdecode

module gpsdecode_tb();
    reg [0:0] clk_i;
    wire [0:0] reset_i; 


endmodule