// testbench for module ssd

module ssd_testbench();

    reg [0:0] clk_i;
    wire [0:0] reset_i;


endmodule