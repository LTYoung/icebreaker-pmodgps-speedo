module speedo
(
    input [0:0] clk_i,
    input [0:0] rst_i,
    output [0:0] o
);  

    assign o = 1'b0;


endmodule